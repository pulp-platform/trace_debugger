// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Author: Robert Balas (balasr@student.ethz.ch)
// Description: Compress instruction traces and filter them


import trdb_pkg::*;

module trace_debugger
    #(parameter APB_ADDR_WIDTH = 32)
    (input logic                clk_i,
     input logic                rst_ni,

     // data from the cpu
     input logic                ivalid_i, //TODO: pipelined valid
     input logic                iexception_i,
     input logic                interrupt_i,
     input logic [CAUSELEN-1:0] cause_i,
     input logic [XLEN-1:0]     tval_i,
     input logic [PRIVLEN-1:0]  priv_i,
     input logic [XLEN-1:0]     iaddr_i,
     input logic [ILEN-1:0]     instr_i,
     input logic                compressed_i,

     APB_BUS.Slave              apb_slave,

     // generated packets, which go the the udma (or somewhere else)
     output logic [XLEN-1:0]    packet_word_o,
     output logic               packet_word_valid_o,
     input logic                stall_i);

    // general control of this module
    // whether this block is enabled at all
    logic                       trace_enable;
    // if we want to trace
    logic                       trace_activated;
    logic                       packet_after_exception;

    logic                       debug_mode;
    logic                       trace_valid;
    logic                       flush_stream;
    logic                       flush_confirm;

    // to register all inputs
    logic                       ivalid_q, ivalid_d;
    logic                       iexception_q, iexception_d;
    logic                       interrupt_q, interrupt_d;
    logic [CAUSELEN-1:0]        cause_q, cause_d;
    // logic [XLEN-1:0]            tval_d, tval_q;
    logic [PRIVLEN-1:0]         priv_q, priv_d;
    logic [XLEN-1:0]            iaddr_q, iaddr_d;
    logic [ILEN-1:0]            instr_q, instr_d;
    logic                       compressed_q, compressed_d;


    // unused variables for a more extensive implementation
    // riscy doesn't have those features
    logic [XLEN-1:0]            lc_tval;
    logic [CONTEXTLEN-1:0]      tc_context;


    // we have three phases, called next cycle (nc), this cycle (tc) and next
    // cycle (nc), based on which we make decision whether we need to emit a
    // packet or not.
    logic [PRIVLEN-1:0]         nc_priv, tc_priv;
    logic                       nc_privchange, tc_privchange;
    logic                       nc_exception, lc_exception;
    logic                       lc_u_discontinuity;
    logic                       tc_first_qualified;
    logic                       tc_is_branch;
    logic                       tc_branch_taken;
    logic                       tc_qualified, lc_qualified, nc_qualified,
                                nc_unqualified;
    logic                       tc_compressed;
    logic [XLEN-1:0]            tc_iaddr, nc_iaddr;
    logic                       lc_exception_sync;
    logic                       lc_interrupt;

    // pass delayed data
    logic [CAUSELEN-1:0]        lc_cause;
    logic                       lc_interupt;

    // registers to hold onto the input data for a few phases, mostly one
    logic                       interrupt0_q, interrupt0_d;
    logic                       interrupt1_q, interrupt1_d;
    logic [CAUSELEN-1:0]        cause0_q, cause0_d;
    logic [CAUSELEN-1:0]        cause1_q, cause1_d;
    logic [PRIVLEN-1:0]         priv0_q, priv0_d;
    logic                       privchange0_q, privchange0_d;
    logic                       exception0_q, exception0_d,
                                exception1_q, exception1_d,
                                exception2_q, exception2_d;
    logic                       u_discontinuity0_q, u_discontinuity0_d,
                                u_discontinuity1_q, u_discontinuity1_d;
    logic                       is_branch0_q, is_branch0_d;
    logic                       compressed0_q, compressed0_d;
    logic [XLEN-1:0]            iaddr0_q, iaddr0_d;
    logic                       qualified0_q, qualified0_d, qualified1_q,
                                qualified1_d;

    // variables for the branch map
    logic                       branch_map_flush;
    logic                       branch_map_full;
    logic                       branch_map_empty;
    logic [30:0]                branch_map;
    logic [4:0]                 branch_map_cnt;

    // variables for the packet generation
    logic                       packet_valid;
    trdb_format_t               packet_format;
    trdb_subformat_t            packet_subformat;

    // generated packet
    logic [PACKET_LEN-1:0]     packet_bits;
    logic [6:0]                packet_len;
    logic                      packet_gen_valid;

    // packet to word
    logic                      packet_is_read;
    logic [XLEN-1:0]           packet_word;
    logic                      packet_word_valid;

    // Holds data from/to advanced peripheral bus
    logic [31:0]               per_rdata;
    logic                      per_ready;
    logic [31:0]               per_wdata;
    logic [APB_ADDR_WIDTH-1:0] per_addr;
    logic                      per_we;
    logic                      per_valid;

    // software dumping: certain writes to the trace debugger are included in
    // the packet stream
    logic [31:0]               sw_word;
    logic                      sw_valid;
    logic                      sw_grant;

    // timer unit
    logic                      timer_rst;
    logic [TIMER_WIDTH-1:0]    tu_time;
    logic                      tu_grant;
    logic                      tu_valid;
    logic                      tu_req;

    // filter unit
    logic                      apply_filters;
    logic                      trace_selected_priv;
    logic [1:0]                trace_which_priv;
    logic                      trace_range;
    logic [XLEN-1:0]           trace_lower_addr;
    logic [XLEN-1:0]           trace_higher_addr;
    logic                      filter_qualified_decision;

    // TODO: send this to reg
    assign timer_rst = '0;

    // to register all inputs
    assign ivalid_d = ivalid_i;
    assign iexception_d = iexception_i;
    assign interrupt_d = interrupt_i;
    assign cause_d  = cause_i;
    assign priv_d = priv_i;
    assign iaddr_d = iaddr_i;
    assign instr_d = instr_i;
    assign compressed_d = compressed_i;

    // whether we do tracing at all
    assign trace_valid = ivalid_q && debug_mode && trace_enable;
    assign debug_mode = priv_q[PRIVLEN-1];

    // TODO: make this configurationr register mapped
    assign packet_after_exception                      = '1;

`ifndef SYNTHESIS
    trace_valid_and_debug: assert property
    (@(posedge clk_i) disable iff (~rst_ni) (trace_enable |-> debug_mode))
        else $info("[TRDB]    @%t: Tracing works only in debug mode",
                   $time);
`endif

    // buffer variables. Certain variables we need to hold up to three cycles
    assign interrupt0_d = interrupt_q;
    assign interrupt1_d = interrupt0_q;
    assign cause0_d = cause_q;
    assign cause1_d = cause0_q;
    assign priv0_d = priv_q;
    assign exception0_d = iexception_q && ivalid_q;
    assign exception1_d = exception0_q;
    assign exception2_d = exception1_q;
    assign compressed0_d = compressed_q;
    assign iaddr0_d = iaddr_q;

    // assign privchange0_d (below)
    // assign u_discontinuity0_d (below)
    // assign is_branch0_d (below)

    assign u_discontinuity1_d = u_discontinuity0_q;
    // TODO: add feature to have selective tracing, add enable with regmap
    assign qualified0_d = trace_enable && filter_qualified_decision; //& ivalid_q
    assign qualified1_d = qualified0_q;

    // Hook phase related variables up to proper register
    assign nc_priv = priv0_d;
    assign tc_priv = priv0_q;
    assign lc_interrupt = interrupt1_q;
    assign lc_cause = cause1_q;
    assign nc_privchange = privchange0_d;
    assign tc_privchange = privchange0_q;
    assign nc_exception = exception0_d;
    assign lc_exception = exception1_q;
    // with that variable we force another packet after an exception packet, so
    // that we don't need to know the vector table entries
    assign lc_exception_sync = exception2_q;
    assign lc_u_discontinuity = u_discontinuity1_q;
    assign tc_is_branch = is_branch0_q;
    assign nc_qualified = qualified0_d;
    assign tc_qualified = qualified0_q;
    assign lc_qualified = qualified1_q;
    assign tc_compressed = compressed0_q;
    assign nc_iaddr = iaddr0_d;
    assign tc_iaddr = iaddr0_q;
    // assign tc_first_qualified (below)
    // assign tc_branch_taken (below)

    // determine if we are allowed to emit packets

    trdb_filter i_trdb_filter
        (.trace_activated_i(trace_activated),
         .apply_filters_i(apply_filters),
         .trace_selected_priv_i(trace_selected_priv),
         .which_priv_i(trace_which_priv),
         .priv_i(priv_d[1:0]),
         .trace_range_i(trace_range),
         .trace_lower_addr_i(trace_lower_addr),
         .trace_higher_addr_i(trace_higher_addr),
         .iaddr_i(iaddr_d),
         .trace_qualified_o(filter_qualified_decision));


    // decide whether a privilege change occured
    always_comb begin
        privchange0_d = (tc_priv != nc_priv) && ivalid_q;
    end

    // decide whether we have a branch instruction
    // beq, bne, blt, bge, bltu, bgeu, p_bneimm, p_beqimm
    always_comb begin: is_branch
        is_branch0_d
            = ((instr_q & MASK_BEQ)      == MATCH_BEQ) ||
              ((instr_q & MASK_BNE)      == MATCH_BNE) ||
              ((instr_q & MASK_BLT)      == MATCH_BLT) ||
              ((instr_q & MASK_BGE)      == MATCH_BGE) ||
              ((instr_q & MASK_BLTU)     == MATCH_BLTU) ||
              ((instr_q & MASK_BGEU)     == MATCH_BGEU) ||
              ((instr_q & MASK_P_BNEIMM) == MATCH_P_BNEIMM) ||
              ((instr_q & MASK_P_BEQIMM) == MATCH_P_BEQIMM);
    end

    // decide whether we have a unpredictable discontinuity
    // jalr, mret, sret, uret
    always_comb begin: is_discontinuity
        u_discontinuity0_d
            = ((instr_q & MASK_JALR) == MATCH_JALR) ||
              ((instr_q & MASK_MRET) == MATCH_MRET) ||
              ((instr_q & MASK_SRET) == MATCH_SRET) ||
              ((instr_q & MASK_URET) == MATCH_URET);
    end

    // figure out whether we are dealing with the first qualified instruction
    always_comb begin: is_qualified
        tc_first_qualified = !lc_qualified && tc_qualified;
    end

    always_comb begin: becomes_unqualified
        nc_unqualified = !nc_qualified;
    end

    // is this branch taken?
    // TODO: change to tc_compressed? 2 :4
    always_comb begin: is_branch_taken
        tc_branch_taken = tc_compressed ?
                          !(tc_iaddr + 2 == nc_iaddr):
                          !(tc_iaddr + 4 == nc_iaddr);
    end

    // update branch map, careful there is a direct combinatorial path
    trdb_branch_map i_trdb_branch_map
        (.clk_i(clk_i),
         .rst_ni(rst_ni),
         .valid_i(tc_is_branch && trace_valid && tc_qualified),
         .branch_taken_i(tc_branch_taken),
         .flush_i(branch_map_flush),
         .map_o(branch_map),
         .branches_o(branch_map_cnt),
         .is_full_o(branch_map_full),
         .is_empty_o(branch_map_empty));

    // decides, by looking at the history of instructions, whether a packet is
    // necessary or not
    trdb_priority i_trdb_priority
        (.clk_i(clk_i),
         .rst_ni(rst_ni),
         // there might be some data stuck in the
         // pipeline if valid never goes high again (e.g.
         // after wfi), but this shouldnt matter
         .valid_i(trace_valid && tc_qualified),
         .lc_exception_i(lc_exception),
         .lc_exception_sync_i(lc_exception_sync && packet_after_exception),

         .tc_first_qualified_i(tc_first_qualified),
         .nc_unqualified_i(nc_unqualified),

         //input logic  tc_unhalted,
         .tc_privchange_i(tc_privchange),
         //input logic resync & branch_map_cnt

         .lc_u_discontinuity_i(lc_u_discontinuity),

         // input logic  resync
         // input logic  branch_map_nonempty,

         //input logic  nc_halt,
         .nc_exception_i(nc_exception),
         .nc_privchange_i(nc_privchange),
         //input logic  nc_qualified,

         .branch_map_full_i(branch_map_full),

         //input logic  tc_context_change,

         .branch_map_empty_i(branch_map_empty),
         .valid_o(packet_valid),
         .packet_format_o(packet_format),
         .packet_subformat_o(packet_subformat));


    // keep track of time for time packets
    trdb_timer
        #(.TIMER_WIDTH(TIMER_WIDTH))
    i_trdb_timer
        (.clk_i(clk_i),
         .rst_ni(rst_ni),
         .manual_rst_i(timer_rst),
         .tu_req_i(tu_req),
         .tu_valid_o(tu_valid),
         .tu_grant_i(tu_grant),
         .trdb_time_o(tu_time));


    // whole packet generation logic
    trdb_packet_emitter i_trdb_packet_emitter
        (.clk_i(clk_i),
         .rst_ni(rst_ni),
         .packet_format_i(packet_format),
         .packet_subformat_i(packet_subformat),
         .valid_i(packet_valid),
         .interrupt_i(lc_interrupt), // get the value of the trapped instr
         .cause_i(lc_cause),
         .tval_i(lc_tval),
         .priv_i(tc_priv),
         .iaddr_i(tc_iaddr),
         .context_i(tc_context),
         .lc_u_discontinuity_i(lc_u_discontinuity),
         .branch_map_i(branch_map),
         .branch_map_cnt_i(branch_map_cnt),
         .branch_map_empty_i(branch_map_empty),
         .branch_map_full_i(branch_map_full),
         .is_branch_i(tc_is_branch),
         .branch_map_flush_o(branch_map_flush),
         .sw_valid_i(sw_valid),
         .sw_word_i(sw_word),
         .sw_grant_o(sw_grant),
         .tu_valid_i(tu_valid),
         .tu_time_i(tu_time),
         .tu_fulltime_i(tu_fulltime),
         .tu_grant_o(tu_grant),
         .packet_bits_o(packet_bits),
         .packet_len_o(packet_len),
         .packet_valid_o(packet_gen_valid),
         .packet_grant_i(packet_is_read));

    trdb_stream_align8 i_trdb_stream_align
        (.clk_i(clk_i),
         .rst_ni(rst_ni),
         .packet_bits_i(packet_bits),
         .packet_len_i(packet_len),
         .valid_i(packet_gen_valid),
         .grant_o(packet_is_read),
         .flush_stream_i(flush_stream),
         .flush_confirm_o(flush_confirm),
         .data_o(packet_word),
         .valid_o(packet_word_valid));

    assign packet_word_o = packet_word;
    assign packet_word_valid_o = packet_word_valid;

    // TODO: assert that we are not dealing with an unsupported instruction
    always_ff @(posedge clk_i, negedge rst_ni) begin
        if(~rst_ni) begin
            ivalid_q           <= '0;
            iexception_q       <= '0;
            interrupt_q        <= '0;
            cause_q            <= '0;
            priv_q             <= '0;
            iaddr_q            <= '0;
            instr_q            <= '0;
            compressed_q       <= '0;

            interrupt0_q       <= '0;
            interrupt1_q       <= '0;
            cause0_q           <= '0;
            cause1_q           <= '0;
            priv0_q            <= 3'h7; //we always start in M-mode
            exception0_q       <= '0;
            exception1_q       <= '0;
            u_discontinuity0_q <= '0;
            u_discontinuity1_q <= '0;
            is_branch0_q       <= '0;
            compressed0_q      <= '0;
            iaddr0_q           <= '0;
            qualified0_q       <= '0;
            qualified1_q       <= '0;
        end else begin
            ivalid_q     <= ivalid_d;
            iexception_q <= iexception_d;
            interrupt_q  <= interrupt_d;
            cause_q      <= cause_d;
            priv_q       <= priv_d;
            iaddr_q      <= iaddr_d;
            instr_q      <= instr_d;
            compressed_q <= compressed_d;

            if(ivalid_q) begin
                interrupt0_q       <= interrupt0_d;
                interrupt1_q       <= interrupt1_d;
                cause0_q           <= cause0_d;
                cause1_q           <= cause1_d;
                priv0_q            <= priv0_d;
                privchange0_q      <= privchange0_d;
                exception0_q       <= exception0_d;
                exception1_q       <= exception1_d;
                exception2_q       <= exception2_d;
                u_discontinuity0_q <= u_discontinuity0_d;
                u_discontinuity1_q <= u_discontinuity1_d;
                is_branch0_q       <= is_branch0_d;
                compressed0_q      <= compressed0_d;
                iaddr0_q           <= iaddr0_d;
                qualified0_q       <= qualified0_d;
                qualified1_q       <= qualified1_d;
            end
        end
    end

    // Connection to the APB. Used to configure the trace debugger. This is just
    // a translation layer.
    trdb_apb_if
        #(.APB_ADDR_WIDTH(APB_ADDR_WIDTH))
    i_trdb_apb_if
        (.paddr(apb_slave.paddr),
         .pwdata(apb_slave.pwdata),
         .pwrite(apb_slave.pwrite),
         .psel(apb_slave.psel),
         .penable(apb_slave.penable),
         .prdata(apb_slave.prdata),
         .pready(apb_slave.pready),
         .pslverr(apb_slave.pslverr),

         .per_rdata_i(per_rdata),
         .per_ready_i(per_ready),
         .per_wdata_o(per_wdata),
         .per_addr_o(per_addr),
         .per_we_o(per_we),
         .per_valid_o(per_valid));

    // Holds configuration data written from the APB and asserts relevant
    // control signals depending on that
    trdb_reg
        #(.APB_ADDR_WIDTH(APB_ADDR_WIDTH))
    i_trdb_reg
        (.clk_i(clk_i),
         .rst_ni(rst_ni),
         .per_rdata_o(per_rdata),
         .per_ready_o(per_ready),
         .per_wdata_i(per_wdata),
         .per_addr_i(per_addr),
         .per_we_i(per_we),
         .per_valid_i(per_valid),
         .flush_stream_o(flush_stream),
         .flush_confirm_i(flush_confirm),
         .trace_enable_o(trace_enable),
         .trace_activated_o(trace_activated),
         .apply_filters_o(apply_filters),
         .trace_selected_priv_o(trace_selected_priv),
         .trace_which_priv_o(trace_which_priv),
         .trace_range_o(trace_range),
         .trace_lower_addr_o(trace_lower_addr),
         .trace_higher_addr_o(trace_higher_addr),
         .sw_word_o(sw_word),
         .sw_valid_o(sw_valid),
         .sw_grant_i(sw_grant),
         .tu_req_o(tu_req));


endmodule // trace_debugger
